///////////////////////////////////////////////////////////////////////////
// Texas A&M University
// CSCE 616 Hardware Design Verification
// Created by  : Prof. Quinn and Saumil Gogri
///////////////////////////////////////////////////////////////////////////

`include "base_test.sv"
`include "simple_random_test.sv"
`include "multiport_sequential_random_test.sv"
`include "corner_test.sv"
`include "random_test.sv"